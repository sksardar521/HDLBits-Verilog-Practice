module top_module( one );

//Insert your code here
    output one;
    assign one = 1'b1;
    

endmodule
